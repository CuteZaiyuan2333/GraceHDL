module test;

     wire a;
    
     wire y;
    
    assign y = a;
    
endmodule
